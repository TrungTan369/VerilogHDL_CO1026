module implement(

    );
    
endmodule
